library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity vector_lien_ke is
  port (
    k_last: in std_logic_vector(15 downto 0) ;
    k1: out std_logic_vector(15 downto 0) ;
    k2: out std_logic_vector(15 downto 0) ;
    k3: out std_logic_vector(15 downto 0) ;
    k4: out std_logic_vector(15 downto 0) ;
    k5: out std_logic_vector(15 downto 0) ;
    k6: out std_logic_vector(15 downto 0) ;
    k7: out std_logic_vector(15 downto 0)
  ) ;
end vector_lien_ke ; 

architecture arch of vector_lien_ke is
    type Row is array ( 0 to 6 ) of integer range 0 to 330 ;
    type VectorTable is array (0 to 330) of Row;
    constant row0: Row := (0, 1 ,2 ,3 ,4 ,5 ,6);
    constant row1: Row := (1, 7 ,8 ,2 ,0 ,6 ,18);
    constant row2: Row := (2, 8 ,9 ,10 ,3 ,0 ,1);
    constant row3: Row := (3, 2 ,10 ,11 ,12 ,4 ,0);
    constant row4: Row := (4, 0 ,3 ,12 ,13 ,14 ,5);
    constant row5: Row := (5, 6 ,0 ,4 ,14 ,15 ,16);
    constant row6: Row := (6, 18 ,1 ,0 ,5 ,16 ,17);
    constant row7: Row := (7, 19 ,20 ,8 ,1 ,18 ,36);
    constant row8: Row := (8, 20 ,21 ,9 ,2 ,1 ,7);
    constant row9: Row := (9, 21 ,22 ,23 ,10 ,2 ,8);
    constant row10: Row := (10, 9 ,23 ,24 ,11 ,3 ,2);
    constant row11: Row := (11, 10 ,24 ,25 ,26 ,12 ,3);
    constant row12: Row := (12, 3 ,11 ,26 ,27 ,13 ,4);
    constant row13: Row := (13, 4 ,12 ,27 ,28 ,29 ,14);
    constant row14: Row := (14, 5 ,4 ,13 ,29 ,30 ,15);
    constant row15: Row := (15, 16 ,5 ,14 ,30 ,31 ,32);
    constant row16: Row := (16, 17 ,6 ,5 ,15 ,32 ,33);
    constant row17: Row := (17, 35 ,18 ,6 ,16 ,33 ,34);
    constant row18: Row := (18, 36 ,7 ,1 ,6 ,17 ,35);
    constant row19: Row := (19, 37 ,38 ,20 ,7 ,36 ,60);
    constant row20: Row := (20, 38 ,39 ,21 ,8 ,7 ,19);
    constant row21: Row := (21, 39 ,40 ,22 ,9 ,8 ,20);
    constant row22: Row := (22, 40 ,41 ,42 ,23 ,9 ,21);
    constant row23: Row := (23, 22 ,42 ,43 ,24 ,10 ,9);
    constant row24: Row := (24, 23 ,43 ,44 ,25 ,11 ,10);
    constant row25: Row := (25, 24 ,44 ,45 ,46 ,26 ,11);
    constant row26: Row := (26, 11 ,25 ,46 ,47 ,27 ,12);
    constant row27: Row := (27, 12 ,26 ,47 ,48 ,28 ,13);
    constant row28: Row := (28, 13 ,27 ,48 ,49 ,50 ,29);
    constant row29: Row := (29, 14 ,13 ,28 ,50 ,51 ,30);
    constant row30: Row := (30, 15 ,14 ,29 ,51 ,52 ,31);
    constant row31: Row := (31, 32 ,15 ,30 ,52 ,53 ,54);
    constant row32: Row := (32, 33 ,16 ,15 ,31 ,54 ,55);
    constant row33: Row := (33, 34 ,17 ,16 ,32 ,55 ,56);
    constant row34: Row := (34, 58 ,35 ,17 ,33 ,56 ,57);
    constant row35: Row := (35, 59 ,36 ,18 ,17 ,34 ,58);
    constant row36: Row := (36, 60 ,19 ,7 ,18 ,35 ,59);
    constant row37: Row := (37, 61 ,62 ,38 ,19 ,60 ,90);
    constant row38: Row := (38, 62 ,63 ,39 ,20 ,19 ,37);
    constant row39: Row := (39, 63 ,64 ,40 ,21 ,20 ,38);
    constant row40: Row := (40, 64 ,65 ,41 ,22 ,21 ,39);
    constant row41: Row := (41, 65 ,66 ,67 ,42 ,22 ,40);
    constant row42: Row := (42, 41 ,67 ,68 ,43 ,23 ,22);
    constant row43: Row := (43, 42 ,68 ,69 ,44 ,24 ,23);
    constant row44: Row := (44, 43 ,69 ,70 ,45 ,25 ,24);
    constant row45: Row := (45, 44 ,70 ,71 ,72 ,46 ,25);
    constant row46: Row := (46, 25 ,45 ,72 ,73 ,47 ,26);
    constant row47: Row := (47, 26 ,46 ,73 ,74 ,48 ,27);
    constant row48: Row := (48, 27 ,47 ,74 ,75 ,49 ,28);
    constant row49: Row := (49, 28 ,48 ,75 ,76 ,77 ,50);
    constant row50: Row := (50, 29 ,28 ,49 ,77 ,78 ,51);
    constant row51: Row := (51, 30 ,29 ,50 ,78 ,79 ,52);
    constant row52: Row := (52, 31 ,30 ,51 ,79 ,80 ,53);
    constant row53: Row := (53, 54 ,31 ,52 ,80 ,81 ,82);
    constant row54: Row := (54, 55 ,32 ,31 ,53 ,82 ,83);
    constant row55: Row := (55, 56 ,33 ,32 ,54 ,83 ,84);
    constant row56: Row := (56, 57 ,34 ,33 ,55 ,84 ,85);
    constant row57: Row := (57, 87 ,58 ,34 ,56 ,85 ,86);
    constant row58: Row := (58, 88 ,59 ,35 ,34 ,57 ,87);
    constant row59: Row := (59, 89 ,60 ,36 ,35 ,58 ,88);
    constant row60: Row := (60, 90 ,37 ,19 ,36 ,59 ,89);
    constant row61: Row := (61, 91 ,92 ,62 ,37 ,90 ,126);
    constant row62: Row := (62, 92 ,93 ,63 ,38 ,37 ,61);
    constant row63: Row := (63, 93 ,94 ,64 ,39 ,38 ,62);
    constant row64: Row := (64, 94 ,95 ,65 ,40 ,39 ,63);
    constant row65: Row := (65, 95 ,96 ,66 ,41 ,40 ,64);
    constant row66: Row := (66, 96 ,97 ,98 ,67 ,41 ,65);
    constant row67: Row := (67, 66 ,98 ,99 ,68 ,42 ,41);
    constant row68: Row := (68, 67 ,99 ,100 ,69 ,43 ,42);
    constant row69: Row := (69, 68 ,100 ,101 ,70 ,44 ,43);
    constant row70: Row := (70, 69 ,101 ,102 ,71 ,45 ,44);
    constant row71: Row := (71, 70 ,102 ,103 ,104 ,72 ,45);
    constant row72: Row := (72, 45 ,71 ,104 ,105 ,73 ,46);
    constant row73: Row := (73, 46 ,72 ,105 ,106 ,74 ,47);
    constant row74: Row := (74, 47 ,73 ,106 ,107 ,75 ,48);
    constant row75: Row := (75, 48 ,74 ,107 ,108 ,76 ,49);
    constant row76: Row := (76, 49 ,75 ,108 ,109 ,110 ,77);
    constant row77: Row := (77, 50 ,49 ,76 ,110 ,111 ,78);
    constant row78: Row := (78, 51 ,50 ,77 ,111 ,112 ,79);
    constant row79: Row := (79, 52 ,51 ,78 ,112 ,113 ,80);
    constant row80: Row := (80, 53 ,52 ,79 ,113 ,114 ,81);
    constant row81: Row := (81, 82 ,53 ,80 ,114 ,115 ,116);
    constant row82: Row := (82, 83 ,54 ,53 ,81 ,116 ,117);
    constant row83: Row := (83, 84 ,55 ,54 ,82 ,117 ,118);
    constant row84: Row := (84, 85 ,56 ,55 ,83 ,118 ,119);
    constant row85: Row := (85, 86 ,57 ,56 ,84 ,119 ,120);
    constant row86: Row := (86, 122 ,87 ,57 ,85 ,120 ,121);
    constant row87: Row := (87, 123 ,88 ,58 ,57 ,86 ,122);
    constant row88: Row := (88, 124 ,89 ,59 ,58 ,87 ,123);
    constant row89: Row := (89, 125 ,90 ,60 ,59 ,88 ,124);
    constant row90: Row := (90, 126 ,61 ,37 ,60 ,89 ,125);
    constant row91: Row := (91, 127 ,128 ,92 ,61 ,126 ,168);
    constant row92: Row := (92, 128 ,129 ,93 ,62 ,61 ,91);
    constant row93: Row := (93, 129 ,130 ,94 ,63 ,62 ,92);
    constant row94: Row := (94, 130 ,131 ,95 ,64 ,63 ,93);
    constant row95: Row := (95, 131 ,132 ,96 ,65 ,64 ,94);
    constant row96: Row := (96, 132 ,133 ,97 ,66 ,65 ,95);
    constant row97: Row := (97, 133 ,134 ,135 ,98 ,66 ,96);
    constant row98: Row := (98, 97 ,135 ,136 ,99 ,67 ,66);
    constant row99: Row := (99, 98 ,136 ,137 ,100 ,68 ,67);
    constant row100: Row := (100, 99 ,137 ,138 ,101 ,69 ,68);
    constant row101: Row := (101, 100 ,138 ,139 ,102 ,70 ,69);
    constant row102: Row := (102, 101 ,139 ,140 ,103 ,71 ,70);
    constant row103: Row := (103, 102 ,140 ,141 ,142 ,104 ,71);
    constant row104: Row := (104, 71 ,103 ,142 ,143 ,105 ,72);
    constant row105: Row := (105, 72 ,104 ,143 ,144 ,106 ,73);
    constant row106: Row := (106, 73 ,105 ,144 ,145 ,107 ,74);
    constant row107: Row := (107, 74 ,106 ,145 ,146 ,108 ,75);
    constant row108: Row := (108, 75 ,107 ,146 ,147 ,109 ,76);
    constant row109: Row := (109, 76 ,108 ,147 ,148 ,149 ,110);
    constant row110: Row := (110, 77 ,76 ,109 ,149 ,150 ,111);
    constant row111: Row := (111, 78 ,77 ,110 ,150 ,151 ,112);
    constant row112: Row := (112, 79 ,78 ,111 ,151 ,152 ,113);
    constant row113: Row := (113, 80 ,79 ,112 ,152 ,153 ,114);
    constant row114: Row := (114, 81 ,80 ,113 ,153 ,154 ,115);
    constant row115: Row := (115, 116 ,81 ,114 ,154 ,155 ,156);
    constant row116: Row := (116, 117 ,82 ,81 ,115 ,156 ,157);
    constant row117: Row := (117, 118 ,83 ,82 ,116 ,157 ,158);
    constant row118: Row := (118, 119 ,84 ,83 ,117 ,158 ,159);
    constant row119: Row := (119, 120 ,85 ,84 ,118 ,159 ,160);
    constant row120: Row := (120, 121 ,86 ,85 ,119 ,160 ,161);
    constant row121: Row := (121, 163 ,122 ,86 ,120 ,161 ,162);
    constant row122: Row := (122, 164 ,123 ,87 ,86 ,121 ,163);
    constant row123: Row := (123, 165 ,124 ,88 ,87 ,122 ,164);
    constant row124: Row := (124, 166 ,125 ,89 ,88 ,123 ,165);
    constant row125: Row := (125, 167 ,126 ,90 ,89 ,124 ,166);
    constant row126: Row := (126, 168 ,91 ,61 ,90 ,125 ,167);
    constant row127: Row := (127, 169 ,170 ,128 ,91 ,168 ,216);
    constant row128: Row := (128, 170 ,171 ,129 ,92 ,91 ,127);
    constant row129: Row := (129, 171 ,172 ,130 ,93 ,92 ,128);
    constant row130: Row := (130, 172 ,173 ,131 ,94 ,93 ,129);
    constant row131: Row := (131, 173 ,174 ,132 ,95 ,94 ,130);
    constant row132: Row := (132, 174 ,175 ,133 ,96 ,95 ,131);
    constant row133: Row := (133, 175 ,176 ,134 ,97 ,96 ,132);
    constant row134: Row := (134, 176 ,177 ,178 ,135 ,97 ,133);
    constant row135: Row := (135, 134 ,178 ,179 ,136 ,98 ,97);
    constant row136: Row := (136, 135 ,179 ,180 ,137 ,99 ,98);
    constant row137: Row := (137, 136 ,180 ,181 ,138 ,100 ,99);
    constant row138: Row := (138, 137 ,181 ,182 ,139 ,101 ,100);
    constant row139: Row := (139, 138 ,182 ,183 ,140 ,102 ,101);
    constant row140: Row := (140, 139 ,183 ,184 ,141 ,103 ,102);
    constant row141: Row := (141, 140 ,184 ,185 ,186 ,142 ,103);
    constant row142: Row := (142, 103 ,141 ,186 ,187 ,143 ,104);
    constant row143: Row := (143, 104 ,142 ,187 ,188 ,144 ,105);
    constant row144: Row := (144, 105 ,143 ,188 ,189 ,145 ,106);
    constant row145: Row := (145, 106 ,144 ,189 ,190 ,146 ,107);
    constant row146: Row := (146, 107 ,145 ,190 ,191 ,147 ,108);
    constant row147: Row := (147, 108 ,146 ,191 ,192 ,148 ,109);
    constant row148: Row := (148, 109 ,147 ,192 ,193 ,194 ,149);
    constant row149: Row := (149, 110 ,109 ,148 ,194 ,195 ,150);
    constant row150: Row := (150, 111 ,110 ,149 ,195 ,196 ,151);
    constant row151: Row := (151, 112 ,111 ,150 ,196 ,197 ,152);
    constant row152: Row := (152, 113 ,112 ,151 ,197 ,198 ,153);
    constant row153: Row := (153, 114 ,113 ,152 ,198 ,199 ,154);
    constant row154: Row := (154, 115 ,114 ,153 ,199 ,200 ,155);
    constant row155: Row := (155, 156 ,115 ,154 ,200 ,201 ,202);
    constant row156: Row := (156, 157 ,116 ,115 ,155 ,202 ,203);
    constant row157: Row := (157, 158 ,117 ,116 ,156 ,203 ,204);
    constant row158: Row := (158, 159 ,118 ,117 ,157 ,204 ,205);
    constant row159: Row := (159, 160 ,119 ,118 ,158 ,205 ,206);
    constant row160: Row := (160, 161 ,120 ,119 ,159 ,206 ,207);
    constant row161: Row := (161, 162 ,121 ,120 ,160 ,207 ,208);
    constant row162: Row := (162, 210 ,163 ,121 ,161 ,208 ,209);
    constant row163: Row := (163, 211 ,164 ,122 ,121 ,162 ,210);
    constant row164: Row := (164, 212 ,165 ,123 ,122 ,163 ,211);
    constant row165: Row := (165, 213 ,166 ,124 ,123 ,164 ,212);
    constant row166: Row := (166, 214 ,167 ,125 ,124 ,165 ,213);
    constant row167: Row := (167, 215 ,168 ,126 ,125 ,166 ,214);
    constant row168: Row := (168, 216 ,127 ,91 ,126 ,167 ,215);
    constant row169: Row := (169, 217 ,218 ,170 ,127 ,216 ,270);
    constant row170: Row := (170, 218 ,219 ,171 ,128 ,127 ,169);
    constant row171: Row := (171, 219 ,220 ,172 ,129 ,128 ,170);
    constant row172: Row := (172, 220 ,221 ,173 ,130 ,129 ,171);
    constant row173: Row := (173, 221 ,222 ,174 ,131 ,130 ,172);
    constant row174: Row := (174, 222 ,223 ,175 ,132 ,131 ,173);
    constant row175: Row := (175, 223 ,224 ,176 ,133 ,132 ,174);
    constant row176: Row := (176, 224 ,225 ,177 ,134 ,133 ,175);
    constant row177: Row := (177, 225 ,226 ,227 ,178 ,134 ,176);
    constant row178: Row := (178, 177 ,227 ,228 ,179 ,135 ,134);
    constant row179: Row := (179, 178 ,228 ,229 ,180 ,136 ,135);
    constant row180: Row := (180, 179 ,229 ,230 ,181 ,137 ,136);
    constant row181: Row := (181, 180 ,230 ,231 ,182 ,138 ,137);
    constant row182: Row := (182, 181 ,231 ,232 ,183 ,139 ,138);
    constant row183: Row := (183, 182 ,232 ,233 ,184 ,140 ,139);
    constant row184: Row := (184, 183 ,233 ,234 ,185 ,141 ,140);
    constant row185: Row := (185, 184 ,234 ,235 ,236 ,186 ,141);
    constant row186: Row := (186, 141 ,185 ,236 ,237 ,187 ,142);
    constant row187: Row := (187, 142 ,186 ,237 ,238 ,188 ,143);
    constant row188: Row := (188, 143 ,187 ,238 ,239 ,189 ,144);
    constant row189: Row := (189, 144 ,188 ,239 ,240 ,190 ,145);
    constant row190: Row := (190, 145 ,189 ,240 ,241 ,191 ,146);
    constant row191: Row := (191, 146 ,190 ,241 ,242 ,192 ,147);
    constant row192: Row := (192, 147 ,191 ,242 ,243 ,193 ,148);
    constant row193: Row := (193, 148 ,192 ,243 ,244 ,245 ,194);
    constant row194: Row := (194, 149 ,148 ,193 ,245 ,246 ,195);
    constant row195: Row := (195, 150 ,149 ,194 ,246 ,247 ,196);
    constant row196: Row := (196, 151 ,150 ,195 ,247 ,248 ,197);
    constant row197: Row := (197, 152 ,151 ,196 ,248 ,249 ,198);
    constant row198: Row := (198, 153 ,152 ,197 ,249 ,250 ,199);
    constant row199: Row := (199, 154 ,153 ,198 ,250 ,251 ,200);
    constant row200: Row := (200, 155 ,154 ,199 ,251 ,252 ,201);
    constant row201: Row := (201, 202 ,155 ,200 ,252 ,253 ,254);
    constant row202: Row := (202, 203 ,156 ,155 ,201 ,254 ,255);
    constant row203: Row := (203, 204 ,157 ,156 ,202 ,255 ,256);
    constant row204: Row := (204, 205 ,158 ,157 ,203 ,256 ,257);
    constant row205: Row := (205, 206 ,159 ,158 ,204 ,257 ,258);
    constant row206: Row := (206, 207 ,160 ,159 ,205 ,258 ,259);
    constant row207: Row := (207, 208 ,161 ,160 ,206 ,259 ,260);
    constant row208: Row := (208, 209 ,162 ,161 ,207 ,260 ,261);
    constant row209: Row := (209, 263 ,210 ,162 ,208 ,261 ,262);
    constant row210: Row := (210, 264 ,211 ,163 ,162 ,209 ,263);
    constant row211: Row := (211, 265 ,212 ,164 ,163 ,210 ,264);
    constant row212: Row := (212, 266 ,213 ,165 ,164 ,211 ,265);
    constant row213: Row := (213, 267 ,214 ,166 ,165 ,212 ,266);
    constant row214: Row := (214, 268 ,215 ,167 ,166 ,213 ,267);
    constant row215: Row := (215, 269 ,216 ,168 ,167 ,214 ,268);
    constant row216: Row := (216, 270 ,169 ,127 ,168 ,215 ,269);
    constant row217: Row := (217, 271 ,272 ,218 ,169 ,270 ,330);
    constant row218: Row := (218, 272 ,273 ,219 ,170 ,169 ,217);
    constant row219: Row := (219, 273 ,274 ,220 ,171 ,170 ,218);
    constant row220: Row := (220, 274 ,275 ,221 ,172 ,171 ,219);
    constant row221: Row := (221, 275 ,276 ,222 ,173 ,172 ,220);
    constant row222: Row := (222, 276 ,277 ,223 ,174 ,173 ,221);
    constant row223: Row := (223, 277 ,278 ,224 ,175 ,174 ,222);
    constant row224: Row := (224, 278 ,279 ,225 ,176 ,175 ,223);
    constant row225: Row := (225, 279 ,280 ,226 ,177 ,176 ,224);
    constant row226: Row := (226, 280 ,281 ,282 ,227 ,177 ,225);
    constant row227: Row := (227, 226 ,282 ,283 ,228 ,178 ,177);
    constant row228: Row := (228, 227 ,283 ,284 ,229 ,179 ,178);
    constant row229: Row := (229, 228 ,284 ,285 ,230 ,180 ,179);
    constant row230: Row := (230, 229 ,285 ,286 ,231 ,181 ,180);
    constant row231: Row := (231, 230 ,286 ,287 ,232 ,182 ,181);
    constant row232: Row := (232, 231 ,287 ,288 ,233 ,183 ,182);
    constant row233: Row := (233, 232 ,288 ,289 ,234 ,184 ,183);
    constant row234: Row := (234, 233 ,289 ,290 ,235 ,185 ,184);
    constant row235: Row := (235, 234 ,290 ,291 ,292 ,236 ,185);
    constant row236: Row := (236, 185 ,235 ,292 ,293 ,237 ,186);
    constant row237: Row := (237, 186 ,236 ,293 ,294 ,238 ,187);
    constant row238: Row := (238, 187 ,237 ,294 ,295 ,239 ,188);
    constant row239: Row := (239, 188 ,238 ,295 ,296 ,240 ,189);
    constant row240: Row := (240, 189 ,239 ,296 ,297 ,241 ,190);
    constant row241: Row := (241, 190 ,240 ,297 ,298 ,242 ,191);
    constant row242: Row := (242, 191 ,241 ,298 ,299 ,243 ,192);
    constant row243: Row := (243, 192 ,242 ,299 ,300 ,244 ,193);
    constant row244: Row := (244, 193 ,243 ,300 ,301 ,302 ,245);
    constant row245: Row := (245, 194 ,193 ,244 ,302 ,303 ,246);
    constant row246: Row := (246, 195 ,194 ,245 ,303 ,304 ,247);
    constant row247: Row := (247, 196 ,195 ,246 ,304 ,305 ,248);
    constant row248: Row := (248, 197 ,196 ,247 ,305 ,306 ,249);
    constant row249: Row := (249, 198 ,197 ,248 ,306 ,307 ,250);
    constant row250: Row := (250, 199 ,198 ,249 ,307 ,308 ,251);
    constant row251: Row := (251, 200 ,199 ,250 ,308 ,309 ,252);
    constant row252: Row := (252, 201 ,200 ,251 ,309 ,310 ,253);
    constant row253: Row := (253, 254 ,201 ,252 ,310 ,311 ,312);
    constant row254: Row := (254, 255 ,202 ,201 ,253 ,312 ,313);
    constant row255: Row := (255, 256 ,203 ,202 ,254 ,313 ,314);
    constant row256: Row := (256, 257 ,204 ,203 ,255 ,314 ,315);
    constant row257: Row := (257, 258 ,205 ,204 ,256 ,315 ,316);
    constant row258: Row := (258, 259 ,206 ,205 ,257 ,316 ,317);
    constant row259: Row := (259, 260 ,207 ,206 ,258 ,317 ,318);
    constant row260: Row := (260, 261 ,208 ,207 ,259 ,318 ,319);
    constant row261: Row := (261, 262 ,209 ,208 ,260 ,319 ,320);
    constant row262: Row := (262, 322 ,263 ,209 ,261 ,320 ,321);
    constant row263: Row := (263, 323 ,264 ,210 ,209 ,262 ,322);
    constant row264: Row := (264, 324 ,265 ,211 ,210 ,263 ,323);
    constant row265: Row := (265, 325 ,266 ,212 ,211 ,264 ,324);
    constant row266: Row := (266, 326 ,267 ,213 ,212 ,265 ,325);
    constant row267: Row := (267, 327 ,268 ,214 ,213 ,266 ,326);
    constant row268: Row := (268, 328 ,269 ,215 ,214 ,267 ,327);
    constant row269: Row := (269, 329 ,270 ,216 ,215 ,268 ,328);
    constant row270: Row := (270, 330 ,217 ,169 ,216 ,269 ,329);
    constant row271: Row := (271, 271 ,217 ,272 ,217 ,330 ,271);
    constant row272: Row := (272, 271 ,217 ,273 ,218 ,217 ,271);
    constant row273: Row := (273, 271 ,217 ,274 ,219 ,218 ,272);
    constant row274: Row := (274, 271 ,217 ,275 ,220 ,219 ,273);
    constant row275: Row := (275, 271 ,217 ,276 ,221 ,220 ,274);
    constant row276: Row := (276, 271 ,217 ,277 ,222 ,221 ,275);
    constant row277: Row := (277, 271 ,217 ,278 ,223 ,222 ,276);
    constant row278: Row := (278, 271 ,217 ,279 ,224 ,223 ,277);
    constant row279: Row := (279, 271 ,217 ,280 ,225 ,224 ,278);
    constant row280: Row := (280, 271 ,217 ,281 ,226 ,225 ,279);
    constant row281: Row := (281, 271 ,281 ,281 ,282 ,226 ,280);
    constant row282: Row := (282, 281 ,282 ,282 ,283 ,227 ,226);
    constant row283: Row := (283, 282 ,283 ,283 ,284 ,228 ,227);
    constant row284: Row := (284, 283 ,284 ,284 ,285 ,229 ,228);
    constant row285: Row := (285, 284 ,285 ,285 ,286 ,230 ,229);
    constant row286: Row := (286, 285 ,286 ,286 ,287 ,231 ,230);
    constant row287: Row := (287, 286 ,287 ,287 ,288 ,232 ,231);
    constant row288: Row := (288, 287 ,288 ,288 ,289 ,233 ,232);
    constant row289: Row := (289, 288 ,289 ,289 ,290 ,234 ,233);
    constant row290: Row := (290, 289 ,290 ,290 ,291 ,235 ,234);
    constant row291: Row := (291, 290 ,291 ,291 ,291 ,292 ,235);
    constant row292: Row := (292, 235 ,291 ,292 ,292 ,293 ,236);
    constant row293: Row := (293, 236 ,292 ,293 ,293 ,294 ,237);
    constant row294: Row := (294, 237 ,293 ,294 ,294 ,295 ,238);
    constant row295: Row := (295, 238 ,294 ,295 ,295 ,296 ,239);
    constant row296: Row := (296, 239 ,295 ,296 ,296 ,297 ,240);
    constant row297: Row := (297, 240 ,296 ,297 ,297 ,298 ,241);
    constant row298: Row := (298, 241 ,297 ,298 ,298 ,299 ,242);
    constant row299: Row := (299, 242 ,298 ,299 ,299 ,300 ,243);
    constant row300: Row := (300, 243 ,299 ,300 ,300 ,301 ,244);
    constant row301: Row := (301, 244 ,300 ,301 ,301 ,301 ,302);
    constant row302: Row := (302, 245 ,244 ,301 ,301 ,301 ,303);
    constant row303: Row := (303, 246 ,245 ,302 ,301 ,301 ,304);
    constant row304: Row := (304, 247 ,246 ,303 ,301 ,301 ,305);
    constant row305: Row := (305, 248 ,247 ,304 ,301 ,301 ,306);
    constant row306: Row := (306, 249 ,248 ,305 ,301 ,301 ,307);
    constant row307: Row := (307, 250 ,249 ,306 ,301 ,301 ,308);
    constant row308: Row := (308, 251 ,250 ,307 ,301 ,301 ,309);
    constant row309: Row := (309, 252 ,251 ,308 ,301 ,301 ,310);
    constant row310: Row := (310, 253 ,252 ,309 ,301 ,301 ,311);
    constant row311: Row := (311, 312 ,253 ,310 ,301 ,311 ,311);
    constant row312: Row := (312, 313 ,254 ,253 ,311 ,312 ,312);
    constant row313: Row := (313, 314 ,255 ,254 ,312 ,313 ,313);
    constant row314: Row := (314, 315 ,256 ,255 ,313 ,314 ,314);
    constant row315: Row := (315, 316 ,257 ,256 ,314 ,315 ,315);
    constant row316: Row := (316, 317 ,258 ,257 ,315 ,316 ,316);
    constant row317: Row := (317, 318 ,259 ,258 ,316 ,317 ,317);
    constant row318: Row := (318, 319 ,260 ,259 ,317 ,318 ,318);
    constant row319: Row := (319, 320 ,261 ,260 ,318 ,319 ,319);
    constant row320: Row := (320, 321 ,262 ,261 ,319 ,320 ,320);
    constant row321: Row := (321, 321 ,322 ,262 ,320 ,321 ,321);
    constant row322: Row := (322, 322 ,323 ,263 ,262 ,321 ,322);
    constant row323: Row := (323, 323 ,324 ,264 ,263 ,322 ,323);
    constant row324: Row := (324, 324 ,325 ,265 ,264 ,323 ,324);
    constant row325: Row := (325, 325 ,326 ,266 ,265 ,324 ,325);
    constant row326: Row := (326, 326 ,327 ,267 ,266 ,325 ,326);
    constant row327: Row := (327, 327 ,328 ,268 ,267 ,326 ,327);
    constant row328: Row := (328, 328 ,329 ,269 ,268 ,327 ,328);
    constant row329: Row := (329, 329 ,330 ,270 ,269 ,328 ,329);
    constant row330: Row := (330, 330 ,271 ,217 ,270 ,329 ,330);
    
    constant Vectors: VectorTable := (
        row0,
        row1,
        row2,
        row3,
        row4,
        row5,
        row6,
        row7,
        row8,
        row9,
        row10,
        row11,
        row12,
        row13,
        row14,
        row15,
        row16,
        row17,
        row18,
        row19,
        row20,
        row21,
        row22,
        row23,
        row24,
        row25,
        row26,
        row27,
        row28,
        row29,
        row30,
        row31,
        row32,
        row33,
        row34,
        row35,
        row36,
        row37,
        row38,
        row39,
        row40,
        row41,
        row42,
        row43,
        row44,
        row45,
        row46,
        row47,
        row48,
        row49,
        row50,
        row51,
        row52,
        row53,
        row54,
        row55,
        row56,
        row57,
        row58,
        row59,
        row60,
        row61,
        row62,
        row63,
        row64,
        row65,
        row66,
        row67,
        row68,
        row69,
        row70,
        row71,
        row72,
        row73,
        row74,
        row75,
        row76,
        row77,
        row78,
        row79,
        row80,
        row81,
        row82,
        row83,
        row84,
        row85,
        row86,
        row87,
        row88,
        row89,
        row90,
        row91,
        row92,
        row93,
        row94,
        row95,
        row96,
        row97,
        row98,
        row99,
        row100,
        row101,
        row102,
        row103,
        row104,
        row105,
        row106,
        row107,
        row108,
        row109,
        row110,
        row111,
        row112,
        row113,
        row114,
        row115,
        row116,
        row117,
        row118,
        row119,
        row120,
        row121,
        row122,
        row123,
        row124,
        row125,
        row126,
        row127,
        row128,
        row129,
        row130,
        row131,
        row132,
        row133,
        row134,
        row135,
        row136,
        row137,
        row138,
        row139,
        row140,
        row141,
        row142,
        row143,
        row144,
        row145,
        row146,
        row147,
        row148,
        row149,
        row150,
        row151,
        row152,
        row153,
        row154,
        row155,
        row156,
        row157,
        row158,
        row159,
        row160,
        row161,
        row162,
        row163,
        row164,
        row165,
        row166,
        row167,
        row168,
        row169,
        row170,
        row171,
        row172,
        row173,
        row174,
        row175,
        row176,
        row177,
        row178,
        row179,
        row180,
        row181,
        row182,
        row183,
        row184,
        row185,
        row186,
        row187,
        row188,
        row189,
        row190,
        row191,
        row192,
        row193,
        row194,
        row195,
        row196,
        row197,
        row198,
        row199,
        row200,
        row201,
        row202,
        row203,
        row204,
        row205,
        row206,
        row207,
        row208,
        row209,
        row210,
        row211,
        row212,
        row213,
        row214,
        row215,
        row216,
        row217,
        row218,
        row219,
        row220,
        row221,
        row222,
        row223,
        row224,
        row225,
        row226,
        row227,
        row228,
        row229,
        row230,
        row231,
        row232,
        row233,
        row234,
        row235,
        row236,
        row237,
        row238,
        row239,
        row240,
        row241,
        row242,
        row243,
        row244,
        row245,
        row246,
        row247,
        row248,
        row249,
        row250,
        row251,
        row252,
        row253,
        row254,
        row255,
        row256,
        row257,
        row258,
        row259,
        row260,
        row261,
        row262,
        row263,
        row264,
        row265,
        row266,
        row267,
        row268,
        row269,
        row270,
        row271,
        row272,
        row273,
        row274,
        row275,
        row276,
        row277,
        row278,
        row279,
        row280,
        row281,
        row282,
        row283,
        row284,
        row285,
        row286,
        row287,
        row288,
        row289,
        row290,
        row291,
        row292,
        row293,
        row294,
        row295,
        row296,
        row297,
        row298,
        row299,
        row300,
        row301,
        row302,
        row303,
        row304,
        row305,
        row306,
        row307,
        row308,
        row309,
        row310,
        row311,
        row312,
        row313,
        row314,
        row315,
        row316,
        row317,
        row318,
        row319,
        row320,
        row321,
        row322,
        row323,
        row324,
        row325,
        row326,
        row327,
        row328,
        row329,
        row330
    );

begin
    identifier : process( k_last )
    variable k: integer range 0 to 330;
    variable j1, j2, j3, j4, j5, j6, j7: integer range 0 to 331;
    variable rowk: Row;
    begin
        k := to_integer(unsigned(k_last));
        rowk := Vectors(k);
        j1 := rowk(0);
        j2 := rowk(1);
        j3 := rowk(2);
        j4 := rowk(3);
        j5 := rowk(4);
        j6 := rowk(5);
        j7 := rowk(6);
        
        k1 <= std_logic_vector(to_unsigned(j1, 16));
        k2 <= std_logic_vector(to_unsigned(j2, 16));
        k3 <= std_logic_vector(to_unsigned(j3, 16));
        k4 <= std_logic_vector(to_unsigned(j4, 16));
        k5 <= std_logic_vector(to_unsigned(j5, 16));
        k6 <= std_logic_vector(to_unsigned(j6, 16));
        k7 <= std_logic_vector(to_unsigned(j7, 16));
    end process ; -- identifier
end architecture ;