library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity StateLevel11 is
  port (
    Vno: in std_logic_vector(15 downto 0) ;

    Van: out std_logic_vector(3 downto 0) ;
    Vbn: out std_logic_vector(3 downto 0) ;
    Vcn: out std_logic_vector(3 downto 0) 
  ) ;
end StateLevel11 ; 

architecture arch of StateLevel11 is
type StateLevels is array (0 to 330) of std_logic_vector(3 downto 0) ;
constant StateA: StateLevels := (
    "0101",
    "0110",
    "0101",
    "0101",
    "0100",
    "0101",
    "0101",
    "0110",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0100",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0101",
    "0110",
    "0110",
    "0111",
    "1000",
    "0111",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0011",
    "0010",
    "0011",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "0111",
    "0111",
    "1000",
    "1000",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1010",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0000",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1001",
    "1001",
    "1001",
    "1001",
    "1000",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0010",
    "0001",
    "0001",
    "0001",
    "0001",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0001",
    "0001",
    "0001",
    "0001",
    "0010",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "1000",
    "1001",
    "1001",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1000",
    "0111",
    "0110",
    "0101",
    "0100",
    "0011",
    "0010",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0010",
    "0011",
    "0100",
    "0101",
    "0110",
    "0111",
    "1000",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010"    
);

constant StateB: StateLevels := (
    "0101",
    "0101",
    "0101",
    "0110",
    "0101",
    "0101",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0110",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0100",
    "0100",
    "0100",
    "0101",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0011",
    "0100",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "0111",
    "1000",
    "0111",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0011",
    "0010",
    "0011",
    "0011",
    "0011",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1010",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0000",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0010",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0001",
    "0010",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "1000",
    "1001",
    "1001",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1001",
    "1001",
    "1001",
    "1001",
    "1000",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0010",
    "0001",
    "0001",
    "0001",
    "0001",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0001",
    "0001",
    "0001",
    "0000",
    "0001",
    "0010",
    "0011",
    "0100",
    "0101",
    "0110",
    "0111",
    "1000",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1000",
    "0111",
    "0110",
    "0101",
    "0100",
    "0011",
    "0010",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000"    
);

constant StateC: StateLevels := (
    "0101",
    "0101",
    "0100",
    "0101",
    "0101",
    "0110",
    "0101",
    "0100",
    "0100",
    "0100",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0110",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0011",
    "0011",
    "0010",
    "0011",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "0111",
    "1000",
    "0111",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0011",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0000",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1010",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0010",
    "0010",
    "0010",
    "0001",
    "0001",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0001",
    "0001",
    "0010",
    "0010",
    "0010",
    "0011",
    "0100",
    "0100",
    "0101",
    "0110",
    "0110",
    "0111",
    "1000",
    "1000",
    "1000",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1001",
    "1001",
    "1000",
    "1000",
    "1000",
    "0111",
    "0110",
    "0110",
    "0101",
    "0100",
    "0100",
    "0011",
    "0001",
    "0001",
    "0001",
    "0001",
    "0001",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0001",
    "0001",
    "0001",
    "0001",
    "0010",
    "0011",
    "0100",
    "0101",
    "0101",
    "0110",
    "0111",
    "1000",
    "1001",
    "1001",
    "1001",
    "1001",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1001",
    "1001",
    "1001",
    "1001",
    "1000",
    "0111",
    "0110",
    "0101",
    "0101",
    "0100",
    "0011",
    "0010",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0000",
    "0001",
    "0010",
    "0011",
    "0100",
    "0101",
    "0110",
    "0111",
    "1000",
    "1001",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1010",
    "1001",
    "1000",
    "0111",
    "0110",
    "0101",
    "0100",
    "0011",
    "0010",
    "0001"    
);


begin
    identifier : process( Vno )
    variable sVn: unsigned(15 downto 0) ;
    begin
        sVn := unsigned(Vno);
        Van <= StateA(to_integer(sVn));
        Vbn <= StateB(to_integer(sVn));
        Vcn <= StateC(to_integer(sVn));
    end process ; -- identifier
    
end architecture ;