library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity sincoslut is

  port (
    theta: in std_logic_vector(12 downto 0) ;

    sinT: out std_logic_vector(15 downto 0) ;
    cosT: out std_logic_vector(15 downto 0)
    );
    
end sincoslut ; 

architecture arch of sincoslut is
    type Sin_table is array ( 0 to 2047 ) of signed(15 downto 0) ;
    constant CsinTable : Sin_table := (
        x"0000",
        x"0019",
        x"0032",
        x"004B",
        x"0064",
        x"007D",
        x"0096",
        x"00AF",
        x"00C9",
        x"00E2",
        x"00FB",
        x"0114",
        x"012D",
        x"0146",
        x"015F",
        x"0178",
        x"0192",
        x"01AB",
        x"01C4",
        x"01DD",
        x"01F6",
        x"020F",
        x"0228",
        x"0242",
        x"025B",
        x"0274",
        x"028D",
        x"02A6",
        x"02BF",
        x"02D8",
        x"02F1",
        x"030B",
        x"0324",
        x"033D",
        x"0356",
        x"036F",
        x"0388",
        x"03A1",
        x"03BA",
        x"03D4",
        x"03ED",
        x"0406",
        x"041F",
        x"0438",
        x"0451",
        x"046A",
        x"0483",
        x"049C",
        x"04B6",
        x"04CF",
        x"04E8",
        x"0501",
        x"051A",
        x"0533",
        x"054C",
        x"0565",
        x"057F",
        x"0598",
        x"05B1",
        x"05CA",
        x"05E3",
        x"05FC",
        x"0615",
        x"062E",
        x"0647",
        x"0660",
        x"067A",
        x"0693",
        x"06AC",
        x"06C5",
        x"06DE",
        x"06F7",
        x"0710",
        x"0729",
        x"0742",
        x"075B",
        x"0775",
        x"078E",
        x"07A7",
        x"07C0",
        x"07D9",
        x"07F2",
        x"080B",
        x"0824",
        x"083D",
        x"0856",
        x"086F",
        x"0888",
        x"08A2",
        x"08BB",
        x"08D4",
        x"08ED",
        x"0906",
        x"091F",
        x"0938",
        x"0951",
        x"096A",
        x"0983",
        x"099C",
        x"09B5",
        x"09CE",
        x"09E7",
        x"0A00",
        x"0A19",
        x"0A33",
        x"0A4C",
        x"0A65",
        x"0A7E",
        x"0A97",
        x"0AB0",
        x"0AC9",
        x"0AE2",
        x"0AFB",
        x"0B14",
        x"0B2D",
        x"0B46",
        x"0B5F",
        x"0B78",
        x"0B91",
        x"0BAA",
        x"0BC3",
        x"0BDC",
        x"0BF5",
        x"0C0E",
        x"0C27",
        x"0C40",
        x"0C59",
        x"0C72",
        x"0C8B",
        x"0CA4",
        x"0CBD",
        x"0CD6",
        x"0CEF",
        x"0D08",
        x"0D21",
        x"0D3A",
        x"0D53",
        x"0D6C",
        x"0D85",
        x"0D9E",
        x"0DB7",
        x"0DD0",
        x"0DE9",
        x"0E02",
        x"0E1B",
        x"0E34",
        x"0E4D",
        x"0E66",
        x"0E7F",
        x"0E98",
        x"0EB1",
        x"0ECA",
        x"0EE3",
        x"0EFC",
        x"0F15",
        x"0F2E",
        x"0F47",
        x"0F60",
        x"0F79",
        x"0F92",
        x"0FAB",
        x"0FC4",
        x"0FDD",
        x"0FF5",
        x"100E",
        x"1027",
        x"1040",
        x"1059",
        x"1072",
        x"108B",
        x"10A4",
        x"10BD",
        x"10D6",
        x"10EF",
        x"1108",
        x"1121",
        x"1139",
        x"1152",
        x"116B",
        x"1184",
        x"119D",
        x"11B6",
        x"11CF",
        x"11E8",
        x"1201",
        x"1219",
        x"1232",
        x"124B",
        x"1264",
        x"127D",
        x"1296",
        x"12AF",
        x"12C8",
        x"12E0",
        x"12F9",
        x"1312",
        x"132B",
        x"1344",
        x"135D",
        x"1376",
        x"138E",
        x"13A7",
        x"13C0",
        x"13D9",
        x"13F2",
        x"140B",
        x"1423",
        x"143C",
        x"1455",
        x"146E",
        x"1487",
        x"149F",
        x"14B8",
        x"14D1",
        x"14EA",
        x"1503",
        x"151B",
        x"1534",
        x"154D",
        x"1566",
        x"157F",
        x"1597",
        x"15B0",
        x"15C9",
        x"15E2",
        x"15FA",
        x"1613",
        x"162C",
        x"1645",
        x"165D",
        x"1676",
        x"168F",
        x"16A8",
        x"16C0",
        x"16D9",
        x"16F2",
        x"170A",
        x"1723",
        x"173C",
        x"1755",
        x"176D",
        x"1786",
        x"179F",
        x"17B7",
        x"17D0",
        x"17E9",
        x"1802",
        x"181A",
        x"1833",
        x"184C",
        x"1864",
        x"187D",
        x"1896",
        x"18AE",
        x"18C7",
        x"18E0",
        x"18F8",
        x"1911",
        x"192A",
        x"1942",
        x"195B",
        x"1973",
        x"198C",
        x"19A5",
        x"19BD",
        x"19D6",
        x"19EF",
        x"1A07",
        x"1A20",
        x"1A38",
        x"1A51",
        x"1A6A",
        x"1A82",
        x"1A9B",
        x"1AB3",
        x"1ACC",
        x"1AE4",
        x"1AFD",
        x"1B16",
        x"1B2E",
        x"1B47",
        x"1B5F",
        x"1B78",
        x"1B90",
        x"1BA9",
        x"1BC1",
        x"1BDA",
        x"1BF2",
        x"1C0B",
        x"1C24",
        x"1C3C",
        x"1C55",
        x"1C6D",
        x"1C86",
        x"1C9E",
        x"1CB7",
        x"1CCF",
        x"1CE8",
        x"1D00",
        x"1D18",
        x"1D31",
        x"1D49",
        x"1D62",
        x"1D7A",
        x"1D93",
        x"1DAB",
        x"1DC4",
        x"1DDC",
        x"1DF5",
        x"1E0D",
        x"1E25",
        x"1E3E",
        x"1E56",
        x"1E6F",
        x"1E87",
        x"1EA0",
        x"1EB8",
        x"1ED0",
        x"1EE9",
        x"1F01",
        x"1F19",
        x"1F32",
        x"1F4A",
        x"1F63",
        x"1F7B",
        x"1F93",
        x"1FAC",
        x"1FC4",
        x"1FDC",
        x"1FF5",
        x"200D",
        x"2025",
        x"203E",
        x"2056",
        x"206E",
        x"2087",
        x"209F",
        x"20B7",
        x"20D0",
        x"20E8",
        x"2100",
        x"2118",
        x"2131",
        x"2149",
        x"2161",
        x"2179",
        x"2192",
        x"21AA",
        x"21C2",
        x"21DA",
        x"21F3",
        x"220B",
        x"2223",
        x"223B",
        x"2254",
        x"226C",
        x"2284",
        x"229C",
        x"22B4",
        x"22CD",
        x"22E5",
        x"22FD",
        x"2315",
        x"232D",
        x"2345",
        x"235E",
        x"2376",
        x"238E",
        x"23A6",
        x"23BE",
        x"23D6",
        x"23EE",
        x"2407",
        x"241F",
        x"2437",
        x"244F",
        x"2467",
        x"247F",
        x"2497",
        x"24AF",
        x"24C7",
        x"24DF",
        x"24F7",
        x"250F",
        x"2528",
        x"2540",
        x"2558",
        x"2570",
        x"2588",
        x"25A0",
        x"25B8",
        x"25D0",
        x"25E8",
        x"2600",
        x"2618",
        x"2630",
        x"2648",
        x"2660",
        x"2678",
        x"2690",
        x"26A8",
        x"26C0",
        x"26D8",
        x"26EF",
        x"2707",
        x"271F",
        x"2737",
        x"274F",
        x"2767",
        x"277F",
        x"2797",
        x"27AF",
        x"27C7",
        x"27DF",
        x"27F6",
        x"280E",
        x"2826",
        x"283E",
        x"2856",
        x"286E",
        x"2886",
        x"289D",
        x"28B5",
        x"28CD",
        x"28E5",
        x"28FD",
        x"2915",
        x"292C",
        x"2944",
        x"295C",
        x"2974",
        x"298B",
        x"29A3",
        x"29BB",
        x"29D3",
        x"29EB",
        x"2A02",
        x"2A1A",
        x"2A32",
        x"2A49",
        x"2A61",
        x"2A79",
        x"2A91",
        x"2AA8",
        x"2AC0",
        x"2AD8",
        x"2AEF",
        x"2B07",
        x"2B1F",
        x"2B36",
        x"2B4E",
        x"2B66",
        x"2B7D",
        x"2B95",
        x"2BAD",
        x"2BC4",
        x"2BDC",
        x"2BF3",
        x"2C0B",
        x"2C23",
        x"2C3A",
        x"2C52",
        x"2C69",
        x"2C81",
        x"2C98",
        x"2CB0",
        x"2CC8",
        x"2CDF",
        x"2CF7",
        x"2D0E",
        x"2D26",
        x"2D3D",
        x"2D55",
        x"2D6C",
        x"2D84",
        x"2D9B",
        x"2DB3",
        x"2DCA",
        x"2DE2",
        x"2DF9",
        x"2E11",
        x"2E28",
        x"2E3F",
        x"2E57",
        x"2E6E",
        x"2E86",
        x"2E9D",
        x"2EB5",
        x"2ECC",
        x"2EE3",
        x"2EFB",
        x"2F12",
        x"2F29",
        x"2F41",
        x"2F58",
        x"2F6F",
        x"2F87",
        x"2F9E",
        x"2FB5",
        x"2FCD",
        x"2FE4",
        x"2FFB",
        x"3013",
        x"302A",
        x"3041",
        x"3059",
        x"3070",
        x"3087",
        x"309E",
        x"30B6",
        x"30CD",
        x"30E4",
        x"30FB",
        x"3112",
        x"312A",
        x"3141",
        x"3158",
        x"316F",
        x"3186",
        x"319E",
        x"31B5",
        x"31CC",
        x"31E3",
        x"31FA",
        x"3211",
        x"3228",
        x"3240",
        x"3257",
        x"326E",
        x"3285",
        x"329C",
        x"32B3",
        x"32CA",
        x"32E1",
        x"32F8",
        x"330F",
        x"3326",
        x"333D",
        x"3354",
        x"336B",
        x"3382",
        x"3399",
        x"33B0",
        x"33C7",
        x"33DE",
        x"33F5",
        x"340C",
        x"3423",
        x"343A",
        x"3451",
        x"3468",
        x"347F",
        x"3496",
        x"34AD",
        x"34C4",
        x"34DB",
        x"34F2",
        x"3508",
        x"351F",
        x"3536",
        x"354D",
        x"3564",
        x"357B",
        x"3592",
        x"35A8",
        x"35BF",
        x"35D6",
        x"35ED",
        x"3604",
        x"361A",
        x"3631",
        x"3648",
        x"365F",
        x"3675",
        x"368C",
        x"36A3",
        x"36BA",
        x"36D0",
        x"36E7",
        x"36FE",
        x"3714",
        x"372B",
        x"3742",
        x"3758",
        x"376F",
        x"3786",
        x"379C",
        x"37B3",
        x"37CA",
        x"37E0",
        x"37F7",
        x"380D",
        x"3824",
        x"383B",
        x"3851",
        x"3868",
        x"387E",
        x"3895",
        x"38AB",
        x"38C2",
        x"38D8",
        x"38EF",
        x"3906",
        x"391C",
        x"3932",
        x"3949",
        x"395F",
        x"3976",
        x"398C",
        x"39A3",
        x"39B9",
        x"39D0",
        x"39E6",
        x"39FD",
        x"3A13",
        x"3A29",
        x"3A40",
        x"3A56",
        x"3A6C",
        x"3A83",
        x"3A99",
        x"3AAF",
        x"3AC6",
        x"3ADC",
        x"3AF2",
        x"3B09",
        x"3B1F",
        x"3B35",
        x"3B4C",
        x"3B62",
        x"3B78",
        x"3B8E",
        x"3BA5",
        x"3BBB",
        x"3BD1",
        x"3BE7",
        x"3BFD",
        x"3C14",
        x"3C2A",
        x"3C40",
        x"3C56",
        x"3C6C",
        x"3C83",
        x"3C99",
        x"3CAF",
        x"3CC5",
        x"3CDB",
        x"3CF1",
        x"3D07",
        x"3D1D",
        x"3D33",
        x"3D49",
        x"3D60",
        x"3D76",
        x"3D8C",
        x"3DA2",
        x"3DB8",
        x"3DCE",
        x"3DE4",
        x"3DFA",
        x"3E10",
        x"3E26",
        x"3E3C",
        x"3E52",
        x"3E68",
        x"3E7D",
        x"3E93",
        x"3EA9",
        x"3EBF",
        x"3ED5",
        x"3EEB",
        x"3F01",
        x"3F17",
        x"3F2D",
        x"3F43",
        x"3F58",
        x"3F6E",
        x"3F84",
        x"3F9A",
        x"3FB0",
        x"3FC5",
        x"3FDB",
        x"3FF1",
        x"4007",
        x"401D",
        x"4032",
        x"4048",
        x"405E",
        x"4073",
        x"4089",
        x"409F",
        x"40B5",
        x"40CA",
        x"40E0",
        x"40F6",
        x"410B",
        x"4121",
        x"4136",
        x"414C",
        x"4162",
        x"4177",
        x"418D",
        x"41A2",
        x"41B8",
        x"41CE",
        x"41E3",
        x"41F9",
        x"420E",
        x"4224",
        x"4239",
        x"424F",
        x"4264",
        x"427A",
        x"428F",
        x"42A5",
        x"42BA",
        x"42D0",
        x"42E5",
        x"42FA",
        x"4310",
        x"4325",
        x"433B",
        x"4350",
        x"4365",
        x"437B",
        x"4390",
        x"43A5",
        x"43BB",
        x"43D0",
        x"43E5",
        x"43FB",
        x"4410",
        x"4425",
        x"443B",
        x"4450",
        x"4465",
        x"447A",
        x"4490",
        x"44A5",
        x"44BA",
        x"44CF",
        x"44E4",
        x"44FA",
        x"450F",
        x"4524",
        x"4539",
        x"454E",
        x"4563",
        x"4578",
        x"458D",
        x"45A3",
        x"45B8",
        x"45CD",
        x"45E2",
        x"45F7",
        x"460C",
        x"4621",
        x"4636",
        x"464B",
        x"4660",
        x"4675",
        x"468A",
        x"469F",
        x"46B4",
        x"46C9",
        x"46DE",
        x"46F3",
        x"4708",
        x"471C",
        x"4731",
        x"4746",
        x"475B",
        x"4770",
        x"4785",
        x"479A",
        x"47AE",
        x"47C3",
        x"47D8",
        x"47ED",
        x"4802",
        x"4816",
        x"482B",
        x"4840",
        x"4855",
        x"4869",
        x"487E",
        x"4893",
        x"48A8",
        x"48BC",
        x"48D1",
        x"48E6",
        x"48FA",
        x"490F",
        x"4923",
        x"4938",
        x"494D",
        x"4961",
        x"4976",
        x"498A",
        x"499F",
        x"49B4",
        x"49C8",
        x"49DD",
        x"49F1",
        x"4A06",
        x"4A1A",
        x"4A2F",
        x"4A43",
        x"4A58",
        x"4A6C",
        x"4A81",
        x"4A95",
        x"4AA9",
        x"4ABE",
        x"4AD2",
        x"4AE7",
        x"4AFB",
        x"4B0F",
        x"4B24",
        x"4B38",
        x"4B4C",
        x"4B61",
        x"4B75",
        x"4B89",
        x"4B9E",
        x"4BB2",
        x"4BC6",
        x"4BDA",
        x"4BEF",
        x"4C03",
        x"4C17",
        x"4C2B",
        x"4C3F",
        x"4C54",
        x"4C68",
        x"4C7C",
        x"4C90",
        x"4CA4",
        x"4CB8",
        x"4CCC",
        x"4CE1",
        x"4CF5",
        x"4D09",
        x"4D1D",
        x"4D31",
        x"4D45",
        x"4D59",
        x"4D6D",
        x"4D81",
        x"4D95",
        x"4DA9",
        x"4DBD",
        x"4DD1",
        x"4DE5",
        x"4DF9",
        x"4E0D",
        x"4E21",
        x"4E34",
        x"4E48",
        x"4E5C",
        x"4E70",
        x"4E84",
        x"4E98",
        x"4EAC",
        x"4EBF",
        x"4ED3",
        x"4EE7",
        x"4EFB",
        x"4F0F",
        x"4F22",
        x"4F36",
        x"4F4A",
        x"4F5E",
        x"4F71",
        x"4F85",
        x"4F99",
        x"4FAC",
        x"4FC0",
        x"4FD4",
        x"4FE7",
        x"4FFB",
        x"500F",
        x"5022",
        x"5036",
        x"5049",
        x"505D",
        x"5070",
        x"5084",
        x"5097",
        x"50AB",
        x"50BF",
        x"50D2",
        x"50E5",
        x"50F9",
        x"510C",
        x"5120",
        x"5133",
        x"5147",
        x"515A",
        x"516E",
        x"5181",
        x"5194",
        x"51A8",
        x"51BB",
        x"51CE",
        x"51E2",
        x"51F5",
        x"5208",
        x"521C",
        x"522F",
        x"5242",
        x"5255",
        x"5269",
        x"527C",
        x"528F",
        x"52A2",
        x"52B5",
        x"52C9",
        x"52DC",
        x"52EF",
        x"5302",
        x"5315",
        x"5328",
        x"533B",
        x"534E",
        x"5362",
        x"5375",
        x"5388",
        x"539B",
        x"53AE",
        x"53C1",
        x"53D4",
        x"53E7",
        x"53FA",
        x"540D",
        x"5420",
        x"5433",
        x"5445",
        x"5458",
        x"546B",
        x"547E",
        x"5491",
        x"54A4",
        x"54B7",
        x"54CA",
        x"54DC",
        x"54EF",
        x"5502",
        x"5515",
        x"5528",
        x"553A",
        x"554D",
        x"5560",
        x"5572",
        x"5585",
        x"5598",
        x"55AB",
        x"55BD",
        x"55D0",
        x"55E3",
        x"55F5",
        x"5608",
        x"561A",
        x"562D",
        x"5640",
        x"5652",
        x"5665",
        x"5677",
        x"568A",
        x"569C",
        x"56AF",
        x"56C1",
        x"56D4",
        x"56E6",
        x"56F9",
        x"570B",
        x"571D",
        x"5730",
        x"5742",
        x"5755",
        x"5767",
        x"5779",
        x"578C",
        x"579E",
        x"57B0",
        x"57C3",
        x"57D5",
        x"57E7",
        x"57F9",
        x"580C",
        x"581E",
        x"5830",
        x"5842",
        x"5855",
        x"5867",
        x"5879",
        x"588B",
        x"589D",
        x"58AF",
        x"58C1",
        x"58D4",
        x"58E6",
        x"58F8",
        x"590A",
        x"591C",
        x"592E",
        x"5940",
        x"5952",
        x"5964",
        x"5976",
        x"5988",
        x"599A",
        x"59AC",
        x"59BE",
        x"59D0",
        x"59E1",
        x"59F3",
        x"5A05",
        x"5A17",
        x"5A29",
        x"5A3B",
        x"5A4D",
        x"5A5E",
        x"5A70",
        x"5A82",
        x"5A94",
        x"5AA5",
        x"5AB7",
        x"5AC9",
        x"5ADB",
        x"5AEC",
        x"5AFE",
        x"5B10",
        x"5B21",
        x"5B33",
        x"5B45",
        x"5B56",
        x"5B68",
        x"5B79",
        x"5B8B",
        x"5B9D",
        x"5BAE",
        x"5BC0",
        x"5BD1",
        x"5BE3",
        x"5BF4",
        x"5C06",
        x"5C17",
        x"5C29",
        x"5C3A",
        x"5C4B",
        x"5C5D",
        x"5C6E",
        x"5C80",
        x"5C91",
        x"5CA2",
        x"5CB4",
        x"5CC5",
        x"5CD6",
        x"5CE8",
        x"5CF9",
        x"5D0A",
        x"5D1B",
        x"5D2D",
        x"5D3E",
        x"5D4F",
        x"5D60",
        x"5D71",
        x"5D83",
        x"5D94",
        x"5DA5",
        x"5DB6",
        x"5DC7",
        x"5DD8",
        x"5DE9",
        x"5DFA",
        x"5E0B",
        x"5E1C",
        x"5E2D",
        x"5E3F",
        x"5E50",
        x"5E60",
        x"5E71",
        x"5E82",
        x"5E93",
        x"5EA4",
        x"5EB5",
        x"5EC6",
        x"5ED7",
        x"5EE8",
        x"5EF9",
        x"5F0A",
        x"5F1A",
        x"5F2B",
        x"5F3C",
        x"5F4D",
        x"5F5E",
        x"5F6E",
        x"5F7F",
        x"5F90",
        x"5FA0",
        x"5FB1",
        x"5FC2",
        x"5FD3",
        x"5FE3",
        x"5FF4",
        x"6004",
        x"6015",
        x"6026",
        x"6036",
        x"6047",
        x"6057",
        x"6068",
        x"6078",
        x"6089",
        x"6099",
        x"60AA",
        x"60BA",
        x"60CB",
        x"60DB",
        x"60EC",
        x"60FC",
        x"610D",
        x"611D",
        x"612D",
        x"613E",
        x"614E",
        x"615E",
        x"616F",
        x"617F",
        x"618F",
        x"619F",
        x"61B0",
        x"61C0",
        x"61D0",
        x"61E0",
        x"61F1",
        x"6201",
        x"6211",
        x"6221",
        x"6231",
        x"6241",
        x"6251",
        x"6261",
        x"6271",
        x"6282",
        x"6292",
        x"62A2",
        x"62B2",
        x"62C2",
        x"62D2",
        x"62E2",
        x"62F2",
        x"6301",
        x"6311",
        x"6321",
        x"6331",
        x"6341",
        x"6351",
        x"6361",
        x"6371",
        x"6380",
        x"6390",
        x"63A0",
        x"63B0",
        x"63C0",
        x"63CF",
        x"63DF",
        x"63EF",
        x"63FE",
        x"640E",
        x"641E",
        x"642D",
        x"643D",
        x"644D",
        x"645C",
        x"646C",
        x"647B",
        x"648B",
        x"649B",
        x"64AA",
        x"64BA",
        x"64C9",
        x"64D9",
        x"64E8",
        x"64F7",
        x"6507",
        x"6516",
        x"6526",
        x"6535",
        x"6545",
        x"6554",
        x"6563",
        x"6573",
        x"6582",
        x"6591",
        x"65A0",
        x"65B0",
        x"65BF",
        x"65CE",
        x"65DD",
        x"65ED",
        x"65FC",
        x"660B",
        x"661A",
        x"6629",
        x"6639",
        x"6648",
        x"6657",
        x"6666",
        x"6675",
        x"6684",
        x"6693",
        x"66A2",
        x"66B1",
        x"66C0",
        x"66CF",
        x"66DE",
        x"66ED",
        x"66FC",
        x"670B",
        x"671A",
        x"6729",
        x"6737",
        x"6746",
        x"6755",
        x"6764",
        x"6773",
        x"6782",
        x"6790",
        x"679F",
        x"67AE",
        x"67BD",
        x"67CB",
        x"67DA",
        x"67E9",
        x"67F7",
        x"6806",
        x"6815",
        x"6823",
        x"6832",
        x"6840",
        x"684F",
        x"685E",
        x"686C",
        x"687B",
        x"6889",
        x"6898",
        x"68A6",
        x"68B5",
        x"68C3",
        x"68D1",
        x"68E0",
        x"68EE",
        x"68FD",
        x"690B",
        x"6919",
        x"6928",
        x"6936",
        x"6944",
        x"6953",
        x"6961",
        x"696F",
        x"697D",
        x"698C",
        x"699A",
        x"69A8",
        x"69B6",
        x"69C4",
        x"69D3",
        x"69E1",
        x"69EF",
        x"69FD",
        x"6A0B",
        x"6A19",
        x"6A27",
        x"6A35",
        x"6A43",
        x"6A51",
        x"6A5F",
        x"6A6D",
        x"6A7B",
        x"6A89",
        x"6A97",
        x"6AA5",
        x"6AB3",
        x"6AC1",
        x"6ACE",
        x"6ADC",
        x"6AEA",
        x"6AF8",
        x"6B06",
        x"6B13",
        x"6B21",
        x"6B2F",
        x"6B3D",
        x"6B4A",
        x"6B58",
        x"6B66",
        x"6B73",
        x"6B81",
        x"6B8F",
        x"6B9C",
        x"6BAA",
        x"6BB8",
        x"6BC5",
        x"6BD3",
        x"6BE0",
        x"6BEE",
        x"6BFB",
        x"6C09",
        x"6C16",
        x"6C24",
        x"6C31",
        x"6C3F",
        x"6C4C",
        x"6C59",
        x"6C67",
        x"6C74",
        x"6C81",
        x"6C8F",
        x"6C9C",
        x"6CA9",
        x"6CB7",
        x"6CC4",
        x"6CD1",
        x"6CDE",
        x"6CEC",
        x"6CF9",
        x"6D06",
        x"6D13",
        x"6D20",
        x"6D2D",
        x"6D3A",
        x"6D48",
        x"6D55",
        x"6D62",
        x"6D6F",
        x"6D7C",
        x"6D89",
        x"6D96",
        x"6DA3",
        x"6DB0",
        x"6DBD",
        x"6DCA",
        x"6DD6",
        x"6DE3",
        x"6DF0",
        x"6DFD",
        x"6E0A",
        x"6E17",
        x"6E24",
        x"6E30",
        x"6E3D",
        x"6E4A",
        x"6E57",
        x"6E63",
        x"6E70",
        x"6E7D",
        x"6E89",
        x"6E96",
        x"6EA3",
        x"6EAF",
        x"6EBC",
        x"6EC9",
        x"6ED5",
        x"6EE2",
        x"6EEE",
        x"6EFB",
        x"6F07",
        x"6F14",
        x"6F20",
        x"6F2D",
        x"6F39",
        x"6F46",
        x"6F52",
        x"6F5F",
        x"6F6B",
        x"6F77",
        x"6F84",
        x"6F90",
        x"6F9C",
        x"6FA9",
        x"6FB5",
        x"6FC1",
        x"6FCD",
        x"6FDA",
        x"6FE6",
        x"6FF2",
        x"6FFE",
        x"700A",
        x"7016",
        x"7023",
        x"702F",
        x"703B",
        x"7047",
        x"7053",
        x"705F",
        x"706B",
        x"7077",
        x"7083",
        x"708F",
        x"709B",
        x"70A7",
        x"70B3",
        x"70BF",
        x"70CB",
        x"70D6",
        x"70E2",
        x"70EE",
        x"70FA",
        x"7106",
        x"7112",
        x"711D",
        x"7129",
        x"7135",
        x"7141",
        x"714C",
        x"7158",
        x"7164",
        x"716F",
        x"717B",
        x"7186",
        x"7192",
        x"719E",
        x"71A9",
        x"71B5",
        x"71C0",
        x"71CC",
        x"71D7",
        x"71E3",
        x"71EE",
        x"71FA",
        x"7205",
        x"7211",
        x"721C",
        x"7227",
        x"7233",
        x"723E",
        x"7249",
        x"7255",
        x"7260",
        x"726B",
        x"7276",
        x"7282",
        x"728D",
        x"7298",
        x"72A3",
        x"72AF",
        x"72BA",
        x"72C5",
        x"72D0",
        x"72DB",
        x"72E6",
        x"72F1",
        x"72FC",
        x"7307",
        x"7312",
        x"731D",
        x"7328",
        x"7333",
        x"733E",
        x"7349",
        x"7354",
        x"735F",
        x"736A",
        x"7375",
        x"737F",
        x"738A",
        x"7395",
        x"73A0",
        x"73AB",
        x"73B5",
        x"73C0",
        x"73CB",
        x"73D6",
        x"73E0",
        x"73EB",
        x"73F6",
        x"7400",
        x"740B",
        x"7415",
        x"7420",
        x"742B",
        x"7435",
        x"7440",
        x"744A",
        x"7455",
        x"745F",
        x"746A",
        x"7474",
        x"747E",
        x"7489",
        x"7493",
        x"749E",
        x"74A8",
        x"74B2",
        x"74BD",
        x"74C7",
        x"74D1",
        x"74DB",
        x"74E6",
        x"74F0",
        x"74FA",
        x"7504",
        x"750F",
        x"7519",
        x"7523",
        x"752D",
        x"7537",
        x"7541",
        x"754B",
        x"7555",
        x"755F",
        x"7569",
        x"7573",
        x"757D",
        x"7587",
        x"7591",
        x"759B",
        x"75A5",
        x"75AF",
        x"75B9",
        x"75C3",
        x"75CC",
        x"75D6",
        x"75E0",
        x"75EA",
        x"75F4",
        x"75FD",
        x"7607",
        x"7611",
        x"761B",
        x"7624",
        x"762E",
        x"7638",
        x"7641",
        x"764B",
        x"7654",
        x"765E",
        x"7668",
        x"7671",
        x"767B",
        x"7684",
        x"768E",
        x"7697",
        x"76A0",
        x"76AA",
        x"76B3",
        x"76BD",
        x"76C6",
        x"76CF",
        x"76D9",
        x"76E2",
        x"76EB",
        x"76F5",
        x"76FE",
        x"7707",
        x"7710",
        x"771A",
        x"7723",
        x"772C",
        x"7735",
        x"773E",
        x"7747",
        x"7751",
        x"775A",
        x"7763",
        x"776C",
        x"7775",
        x"777E",
        x"7787",
        x"7790",
        x"7799",
        x"77A2",
        x"77AB",
        x"77B4",
        x"77BC",
        x"77C5",
        x"77CE",
        x"77D7",
        x"77E0",
        x"77E9",
        x"77F1",
        x"77FA",
        x"7803",
        x"780C",
        x"7814",
        x"781D",
        x"7826",
        x"782E",
        x"7837",
        x"7840",
        x"7848",
        x"7851",
        x"7859",
        x"7862",
        x"786B",
        x"7873",
        x"787C",
        x"7884",
        x"788C",
        x"7895",
        x"789D",
        x"78A6",
        x"78AE",
        x"78B6",
        x"78BF",
        x"78C7",
        x"78CF",
        x"78D8",
        x"78E0",
        x"78E8",
        x"78F1",
        x"78F9",
        x"7901",
        x"7909",
        x"7911",
        x"7919",
        x"7922",
        x"792A",
        x"7932",
        x"793A",
        x"7942",
        x"794A",
        x"7952",
        x"795A",
        x"7962",
        x"796A",
        x"7972",
        x"797A",
        x"7982",
        x"798A",
        x"7992",
        x"7999",
        x"79A1",
        x"79A9",
        x"79B1",
        x"79B9",
        x"79C0",
        x"79C8",
        x"79D0",
        x"79D8",
        x"79DF",
        x"79E7",
        x"79EF",
        x"79F6",
        x"79FE",
        x"7A05",
        x"7A0D",
        x"7A15",
        x"7A1C",
        x"7A24",
        x"7A2B",
        x"7A33",
        x"7A3A",
        x"7A42",
        x"7A49",
        x"7A50",
        x"7A58",
        x"7A5F",
        x"7A67",
        x"7A6E",
        x"7A75",
        x"7A7D",
        x"7A84",
        x"7A8B",
        x"7A92",
        x"7A9A",
        x"7AA1",
        x"7AA8",
        x"7AAF",
        x"7AB6",
        x"7ABD",
        x"7AC5",
        x"7ACC",
        x"7AD3",
        x"7ADA",
        x"7AE1",
        x"7AE8",
        x"7AEF",
        x"7AF6",
        x"7AFD",
        x"7B04",
        x"7B0B",
        x"7B12",
        x"7B19",
        x"7B1F",
        x"7B26",
        x"7B2D",
        x"7B34",
        x"7B3B",
        x"7B42",
        x"7B48",
        x"7B4F",
        x"7B56",
        x"7B5D",
        x"7B63",
        x"7B6A",
        x"7B71",
        x"7B77",
        x"7B7E",
        x"7B84",
        x"7B8B",
        x"7B92",
        x"7B98",
        x"7B9F",
        x"7BA5",
        x"7BAC",
        x"7BB2",
        x"7BB9",
        x"7BBF",
        x"7BC5",
        x"7BCC",
        x"7BD2",
        x"7BD9",
        x"7BDF",
        x"7BE5",
        x"7BEB",
        x"7BF2",
        x"7BF8",
        x"7BFE",
        x"7C05",
        x"7C0B",
        x"7C11",
        x"7C17",
        x"7C1D",
        x"7C23",
        x"7C29",
        x"7C30",
        x"7C36",
        x"7C3C",
        x"7C42",
        x"7C48",
        x"7C4E",
        x"7C54",
        x"7C5A",
        x"7C60",
        x"7C66",
        x"7C6C",
        x"7C71",
        x"7C77",
        x"7C7D",
        x"7C83",
        x"7C89",
        x"7C8F",
        x"7C94",
        x"7C9A",
        x"7CA0",
        x"7CA6",
        x"7CAB",
        x"7CB1",
        x"7CB7",
        x"7CBC",
        x"7CC2",
        x"7CC8",
        x"7CCD",
        x"7CD3",
        x"7CD8",
        x"7CDE",
        x"7CE3",
        x"7CE9",
        x"7CEE",
        x"7CF4",
        x"7CF9",
        x"7CFF",
        x"7D04",
        x"7D09",
        x"7D0F",
        x"7D14",
        x"7D19",
        x"7D1F",
        x"7D24",
        x"7D29",
        x"7D2F",
        x"7D34",
        x"7D39",
        x"7D3E",
        x"7D43",
        x"7D49",
        x"7D4E",
        x"7D53",
        x"7D58",
        x"7D5D",
        x"7D62",
        x"7D67",
        x"7D6C",
        x"7D71",
        x"7D76",
        x"7D7B",
        x"7D80",
        x"7D85",
        x"7D8A",
        x"7D8F",
        x"7D94",
        x"7D98",
        x"7D9D",
        x"7DA2",
        x"7DA7",
        x"7DAC",
        x"7DB0",
        x"7DB5",
        x"7DBA",
        x"7DBF",
        x"7DC3",
        x"7DC8",
        x"7DCD",
        x"7DD1",
        x"7DD6",
        x"7DDA",
        x"7DDF",
        x"7DE4",
        x"7DE8",
        x"7DED",
        x"7DF1",
        x"7DF6",
        x"7DFA",
        x"7DFF",
        x"7E03",
        x"7E07",
        x"7E0C",
        x"7E10",
        x"7E14",
        x"7E19",
        x"7E1D",
        x"7E21",
        x"7E26",
        x"7E2A",
        x"7E2E",
        x"7E32",
        x"7E37",
        x"7E3B",
        x"7E3F",
        x"7E43",
        x"7E47",
        x"7E4B",
        x"7E4F",
        x"7E53",
        x"7E57",
        x"7E5B",
        x"7E5F",
        x"7E63",
        x"7E67",
        x"7E6B",
        x"7E6F",
        x"7E73",
        x"7E77",
        x"7E7B",
        x"7E7F",
        x"7E83",
        x"7E86",
        x"7E8A",
        x"7E8E",
        x"7E92",
        x"7E95",
        x"7E99",
        x"7E9D",
        x"7EA1",
        x"7EA4",
        x"7EA8",
        x"7EAB",
        x"7EAF",
        x"7EB3",
        x"7EB6",
        x"7EBA",
        x"7EBD",
        x"7EC1",
        x"7EC4",
        x"7EC8",
        x"7ECB",
        x"7ECF",
        x"7ED2",
        x"7ED5",
        x"7ED9",
        x"7EDC",
        x"7EDF",
        x"7EE3",
        x"7EE6",
        x"7EE9",
        x"7EED",
        x"7EF0",
        x"7EF3",
        x"7EF6",
        x"7EF9",
        x"7EFD",
        x"7F00",
        x"7F03",
        x"7F06",
        x"7F09",
        x"7F0C",
        x"7F0F",
        x"7F12",
        x"7F15",
        x"7F18",
        x"7F1B",
        x"7F1E",
        x"7F21",
        x"7F24",
        x"7F27",
        x"7F2A",
        x"7F2D",
        x"7F2F",
        x"7F32",
        x"7F35",
        x"7F38",
        x"7F3B",
        x"7F3D",
        x"7F40",
        x"7F43",
        x"7F45",
        x"7F48",
        x"7F4B",
        x"7F4D",
        x"7F50",
        x"7F53",
        x"7F55",
        x"7F58",
        x"7F5A",
        x"7F5D",
        x"7F5F",
        x"7F62",
        x"7F64",
        x"7F67",
        x"7F69",
        x"7F6B",
        x"7F6E",
        x"7F70",
        x"7F72",
        x"7F75",
        x"7F77",
        x"7F79",
        x"7F7C",
        x"7F7E",
        x"7F80",
        x"7F82",
        x"7F85",
        x"7F87",
        x"7F89",
        x"7F8B",
        x"7F8D",
        x"7F8F",
        x"7F91",
        x"7F93",
        x"7F95",
        x"7F97",
        x"7F99",
        x"7F9B",
        x"7F9D",
        x"7F9F",
        x"7FA1",
        x"7FA3",
        x"7FA5",
        x"7FA7",
        x"7FA9",
        x"7FAA",
        x"7FAC",
        x"7FAE",
        x"7FB0",
        x"7FB1",
        x"7FB3",
        x"7FB5",
        x"7FB7",
        x"7FB8",
        x"7FBA",
        x"7FBC",
        x"7FBD",
        x"7FBF",
        x"7FC0",
        x"7FC2",
        x"7FC3",
        x"7FC5",
        x"7FC6",
        x"7FC8",
        x"7FC9",
        x"7FCB",
        x"7FCC",
        x"7FCE",
        x"7FCF",
        x"7FD0",
        x"7FD2",
        x"7FD3",
        x"7FD4",
        x"7FD6",
        x"7FD7",
        x"7FD8",
        x"7FD9",
        x"7FDA",
        x"7FDC",
        x"7FDD",
        x"7FDE",
        x"7FDF",
        x"7FE0",
        x"7FE1",
        x"7FE2",
        x"7FE3",
        x"7FE4",
        x"7FE5",
        x"7FE6",
        x"7FE7",
        x"7FE8",
        x"7FE9",
        x"7FEA",
        x"7FEB",
        x"7FEC",
        x"7FED",
        x"7FEE",
        x"7FEE",
        x"7FEF",
        x"7FF0",
        x"7FF1",
        x"7FF2",
        x"7FF2",
        x"7FF3",
        x"7FF4",
        x"7FF4",
        x"7FF5",
        x"7FF6",
        x"7FF6",
        x"7FF7",
        x"7FF7",
        x"7FF8",
        x"7FF8",
        x"7FF9",
        x"7FF9",
        x"7FFA",
        x"7FFA",
        x"7FFB",
        x"7FFB",
        x"7FFC",
        x"7FFC",
        x"7FFC",
        x"7FFD",
        x"7FFD",
        x"7FFD",
        x"7FFE",
        x"7FFE",
        x"7FFE",
        x"7FFE",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF",
        x"7FFF"
        
    );

begin
   
    sin_pro : process( theta )
    variable tLookup: unsigned(10 downto 0) ;
    variable amTlookup: unsigned(10 downto 0) ;
    variable sin1, sin2: signed(15 downto 0) ;
    variable t1, t2: integer range 0 to 2047;
    variable sinX, cosX: signed(15 downto 0) ;
    begin
        tLookup := unsigned(theta(10 downto 0));
        amTlookup := 0 - tLookup;

        t1 := to_integer(tLookup);
        t2 := to_integer(amTlookup);

        sin1 := CsinTable(t1);
        sin2 := CsinTable(t2);

        if (tLookup = 0) then
            case( theta(12 downto 11) ) is
        
                when "00" =>
                    sinX := (others => '0');
                    cosX := x"7fff";
                when "01" =>
                    sinX := x"7fff";
                    cosX := (others => '0');
                when "10" =>
                    sinX := (others => '0');
                    cosX := x"8000";
                when "11" =>
                    sinX := x"8000";
                    cosX := (others => '0');
                when others => null;
            
            end case ;
        else
            case( theta(12 downto 11) ) is
        
                when "00" =>
                    sinX := sin1;
                    cosX := sin2;
                when "01" =>
                    sinX := sin2;
                    cosX := 0 - sin1;
                when "10" =>
                    sinX := 0 - sin1;
                    cosX := 0 - sin2;
                when "11" =>
                    sinX := 0 - sin2;
                    cosX := sin1;
                when others => null;
            
            end case ;
        end if ;

        sinT <= std_logic_vector(sinX);
        cost <= std_logic_vector(cosX);
        
    end process ; -- sin_pro

end architecture ;